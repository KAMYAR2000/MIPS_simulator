module Adder(input [15:0] in, pluser, output [15:0] out);
    assign out = in + pluser;
endmodule

////////&