module Jumper(input [15:0] pc, input [11:0] adress, output [15:0] pc_out);
    assign pc_out = {pc[15:13], adress , 1'b0};
endmodule
/////////////////&